
module test2(a,b,c,d,out);
input wire a;
input wire b;
input wire c;
input wire d;
output reg [15:0] out;
always@(*)begin
  case({a,b,c,d})
  4'b0000:out = 16'b0000_0000_0000_0001;
  4'b0001:out = 16'b0000_0000_0000_0010;
  4'b0010:out = 16'b0000_0000_0000_0100;
  4'b0011:out = 16'b0000_0000_0000_1000;
  4'b0100:out = 16'b0000_0000_0001_0000;
  4'b0101:out = 16'b0000_0000_0010_0000;
  4'b0110:out = 16'b0000_0000_0100_0000;
  4'b0111:out = 16'b0000_0000_1000_0000;
  4'b1000:out = 16'b0000_0001_0000_0000;
  4'b1001:out = 16'b0000_0010_0000_0000;
  4'b1010:out = 16'b0000_0100_0000_0000;
  4'b1011:out = 16'b0000_1000_0000_0000;
  4'b1100:out = 16'b0001_0000_0000_0000;
  4'b1101:out = 16'b0010_0000_0000_0000;
  4'b1110:out = 16'b0100_0000_0000_0000;
  4'b1111:out = 16'b1000_0000_0000_0000;
  endcase
  end
endmodule
